library verilog;
use verilog.vl_types.all;
entity Tb_RhythmGame is
end Tb_RhythmGame;
